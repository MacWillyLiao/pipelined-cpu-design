module control_single( opcode, Funct, NOP, RegDst, ALUSrc, MemtoReg, RegWrite, 
					             MemRead, MemWrite, Branch, Jump, ALUOp, JumpR);
    input[5:0] opcode, Funct;
    input NOP ;
    output RegDst, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, Jump, JumpR;
    output[1:0] ALUOp;
    reg RegDst, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, Jump, JumpR;
    reg[1:0] ALUOp;

    parameter R_FORMAT = 6'd0;
    parameter LW = 6'd35;
    parameter SW = 6'd43;
    parameter BEQ = 6'd4;
	  parameter J = 6'd2;
	  parameter ANDI = 6'd12;

    always @( opcode or Funct ) begin
        case ( opcode )
          R_FORMAT : 
          if ( Funct == 6'd8 ) begin
              RegDst = 1'bx; ALUSrc = 1'bx; MemtoReg = 1'bx; RegWrite = 1'b0; MemRead = 1'b0; 
              MemWrite = 1'b0; Branch = 1'b1; Jump = 1'b1; ALUOp = 2'b10; JumpR = 1'b1;
          end else if ( NOP ) begin
              RegDst = 1'b0; ALUSrc = 1'b0; MemtoReg = 1'b0; RegWrite = 1'b0; MemRead = 1'b0; 
              MemWrite = 1'b0; Branch = 1'b0; Jump = 1'b0; ALUOp = 2'b00; JumpR = 1'b0;
          end else begin
				      RegDst = 1'b1; ALUSrc = 1'b0; MemtoReg = 1'b0; RegWrite = 1'b1; MemRead = 1'b0; 
				      MemWrite = 1'b0; Branch = 1'b0; Jump = 1'b0; ALUOp = 2'b10; JumpR = 1'b0;
          end
          LW :
          begin
				RegDst = 1'b0; ALUSrc = 1'b1; MemtoReg = 1'b1; RegWrite = 1'b1; MemRead = 1'b1; 
				MemWrite = 1'b0; Branch = 1'b0; Jump = 1'b0; ALUOp = 2'b00; JumpR = 1'b0;
          end
          SW :
          begin
				RegDst = 1'bx; ALUSrc = 1'b1; MemtoReg = 1'bx; RegWrite = 1'b0; MemRead = 1'b0; 
				MemWrite = 1'b1; Branch = 1'b0; Jump = 1'b0; ALUOp = 2'b00; JumpR = 1'b0;
          end
          BEQ :
          begin
				RegDst = 1'bx; ALUSrc = 1'b0; MemtoReg = 1'bx; RegWrite = 1'b0; MemRead = 1'b0; 
				MemWrite = 1'b0; Branch = 1'b1; Jump = 1'b0; ALUOp = 2'b01; JumpR = 1'b0;
          end
		      J :
		      begin
				RegDst = 1'bx; ALUSrc = 1'b0; MemtoReg = 1'bx; RegWrite = 1'b0; MemRead = 1'b0; 
				MemWrite = 1'b0; Branch = 1'b1; Jump = 1'b1; ALUOp = 2'b01; JumpR = 1'b0;
		      end
		      ANDI :
		      begin
		    RegDst = 1'b0; ALUSrc = 1'b1; MemtoReg = 1'b0; RegWrite = 1'b1; MemRead = 1'b0; 
        MemWrite = 1'b0; Branch = 1'b0; Jump = 1'b0; ALUOp = 2'b11; JumpR = 1'b0;
		      end
          default
          begin
				$display("control_single unimplemented opcode %d", opcode);
				RegDst=1'bx; ALUSrc=1'bx; MemtoReg=1'bx; RegWrite=1'bx; MemRead=1'bx; 
				MemWrite=1'bx; Branch=1'bx; Jump = 1'bx; ALUOp = 2'bxx; JumpR = 1'bx;
          end
        endcase
    end
endmodule

